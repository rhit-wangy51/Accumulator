module mux1b1(
	input [0:0] A,
	input [0:0] B,
	input [0:0] OP,
	output reg [0:0] Out
);


always begin
	if(OP==1'b0)
		Out <= A; 
	else
		Out <= B;
end

endmodule
